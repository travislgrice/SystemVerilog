
`timescale 1ns / 1ps

/* The module is the basic building block for designs. */
module Testbench(logic clock);
    localparam default_opcode = 5'b11010;

    //////////////////////////////////////////////////////////////////////////////
    /* Modules can contain hierarchies of other modules...                      */
    //////////////////////////////////////////////////////////////////////////////
    /*  */
    bit unsigned [4:0] opcode;
    bit unsigned [15:5] address;
    string debug_msg;
    bit error;
    
    module Adapter();
        module Controller();
        endmodule: Controller
        module Encoder();
            module Multiplexer;
            endmodule: Multiplexer
        endmodule: Encoder
    endmodule: Adapter
    
    ///////////////
    /*... nets.. */
    ///////////////
    wire [9:0] primary_connection;
    reg a, b, c;
    
    /*... variables... */
    logic unsigned [15:0] instruction;
    integer mode;
    Adapter adapter();
    
    //////////////////////////////////
    /*... subroutine declarations.. */
    //////////////////////////////////
    
    ///////////////////////////////////////////////////////////////////////
    /*... and procedural statements within always and initial procedures.*/
    ///////////////////////////////////////////////////////////////////////
    initial begin
        opcode = default_opcode;
        debug_msg = "No error discovered.";
        error = 1'b0;
        // encapsulate instruction within opcode and mode
        instruction = {opcode, address};
        
    end
    
    initial begin
        debug_msg = "Starting simulation.";
        $display(debug_msg);
    end
    
    final begin
        debug_msg = "Ending simulation.";
        $display(debug_msg);
    end
   
    always @(posedge clock) begin
        if (instruction == 16'h00) begin
            reset();
        end else begin
            address++;
        end
    end
    
    task reset();
        opcode = default_opcode;
        address = 11'h000;
        debug_msg = "System has been reset";
        error = 1'b1;
        #100;
        error = 1'b0;
        debug_msg = "No error discovered.";
    endtask: reset
    //////////////////////////////////////////////////////////////////////////////
    /* However,  for  the  testbench, the emphasis is not in the hardware-level */
    /* details such  as wires,  structural heirarchy, and interconnects, but in */
    /* modeling the complete  environment  in  which  a design is verified. The */
    /* environment  must  be properly initialized  and  synchronized,  avoiding */
    /* races  between  the design and the testbench, automating the generations */
    /* of input stimuli, and  reusing existing models and other infrastructure. */
    /* See                 notes                 on                 "Programs". */
    //////////////////////////////////////////////////////////////////////////////
    
endmodule

////////////////////////////////////////////////////////////////////////////////
/* The program  construct  serves  as a  clear separator  between design  and */
/* testbench,  and,  more  importantly,  it  specifies  specialized execution */
/* semantics in the reactive region set  for all elements declared within the */
/* program. Together with clocking blocks, the program construct provides for */
/* race-free interaction  between the design  and the testbench  and  enables */
/* cycle-             and             transaction-level         abstractions. */
////////////////////////////////////////////////////////////////////////////////
program First_Program;

    /* A typical program contains type and data declarations... */
    class SGL_Descriptor;
    endclass: SGL_Descriptor
    
    class NVMe_Instruction;
        typedef class Data_Pointer;
        Data_Pointer data_pointer;
        class Data_Pointer;
            // Class items go here.
        endclass: Data_Pointer
    endclass: NVMe_Instruction
    SGL_Descriptor data_block_descriptor = new;
    
    ////////////////////////////////////////////////////////////////////////////////
    /* program_nonansi_header ::=                                                 */
    /*     {attribute_instance}program[lifetime]program_identifier                */
    /*         {package_import_declaration}[parameter_port_list][list_of_port_de] */
    ////////////////////////////////////////////////////////////////////////////////

endprogram: First_Program

package data_package;
endpackage: data_package

(* concurrent *)
program automatic data_process
import data_package::*;
#(time time_slice = 10ms)(input integer data_in, output integer data_out);
    timeunit 1ms;
    timeprecision 100ns;
    // program items go here.
endprogram: data_process

///////////////////////////////////////////////////////////////////////////////////
/* These are a couple of examples (more or less) from the IEEE 1800 specification*/
///////////////////////////////////////////////////////////////////////////////////
program test(input clk, input [16:1] addr, inout [7:0] data);
    initial begin
        // some initializations go here
    end
endprogram: test

program test2(interface device_ifc);
    initial begin
        // some initializations go here
    end
endprogram: test2
